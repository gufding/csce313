// nios_system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module nios_system (
		input  wire        clk_clk,                           //                         clk.clk
		output wire [12:0] new_sdram_controller_0_wire_addr,  // new_sdram_controller_0_wire.addr
		output wire [1:0]  new_sdram_controller_0_wire_ba,    //                            .ba
		output wire        new_sdram_controller_0_wire_cas_n, //                            .cas_n
		output wire        new_sdram_controller_0_wire_cke,   //                            .cke
		output wire        new_sdram_controller_0_wire_cs_n,  //                            .cs_n
		inout  wire [31:0] new_sdram_controller_0_wire_dq,    //                            .dq
		output wire [3:0]  new_sdram_controller_0_wire_dqm,   //                            .dqm
		output wire        new_sdram_controller_0_wire_ras_n, //                            .ras_n
		output wire        new_sdram_controller_0_wire_we_n,  //                            .we_n
		input  wire        reset_reset_n,                     //                       reset.reset_n
		output wire        sdram_clk_clk,                     //                   sdram_clk.clk
		inout  wire [15:0] sram_DQ,                           //                        sram.DQ
		output wire [19:0] sram_ADDR,                         //                            .ADDR
		output wire        sram_LB_N,                         //                            .LB_N
		output wire        sram_UB_N,                         //                            .UB_N
		output wire        sram_CE_N,                         //                            .CE_N
		output wire        sram_OE_N,                         //                            .OE_N
		output wire        sram_WE_N,                         //                            .WE_N
		output wire        vga_CLK,                           //                         vga.CLK
		output wire        vga_HS,                            //                            .HS
		output wire        vga_VS,                            //                            .VS
		output wire        vga_BLANK,                         //                            .BLANK
		output wire        vga_SYNC,                          //                            .SYNC
		output wire [7:0]  vga_R,                             //                            .R
		output wire [7:0]  vga_G,                             //                            .G
		output wire [7:0]  vga_B                              //                            .B
	);

	wire         video_alpha_blender_0_avalon_blended_source_valid;                                        // video_alpha_blender_0:output_valid -> video_dual_clock_buffer_0:stream_in_valid
	wire  [29:0] video_alpha_blender_0_avalon_blended_source_data;                                         // video_alpha_blender_0:output_data -> video_dual_clock_buffer_0:stream_in_data
	wire         video_alpha_blender_0_avalon_blended_source_ready;                                        // video_dual_clock_buffer_0:stream_in_ready -> video_alpha_blender_0:output_ready
	wire         video_alpha_blender_0_avalon_blended_source_startofpacket;                                // video_alpha_blender_0:output_startofpacket -> video_dual_clock_buffer_0:stream_in_startofpacket
	wire         video_alpha_blender_0_avalon_blended_source_endofpacket;                                  // video_alpha_blender_0:output_endofpacket -> video_dual_clock_buffer_0:stream_in_endofpacket
	wire         video_character_buffer_with_dma_0_avalon_char_source_valid;                               // video_character_buffer_with_dma_0:stream_valid -> video_alpha_blender_0:foreground_valid
	wire  [39:0] video_character_buffer_with_dma_0_avalon_char_source_data;                                // video_character_buffer_with_dma_0:stream_data -> video_alpha_blender_0:foreground_data
	wire         video_character_buffer_with_dma_0_avalon_char_source_ready;                               // video_alpha_blender_0:foreground_ready -> video_character_buffer_with_dma_0:stream_ready
	wire         video_character_buffer_with_dma_0_avalon_char_source_startofpacket;                       // video_character_buffer_with_dma_0:stream_startofpacket -> video_alpha_blender_0:foreground_startofpacket
	wire         video_character_buffer_with_dma_0_avalon_char_source_endofpacket;                         // video_character_buffer_with_dma_0:stream_endofpacket -> video_alpha_blender_0:foreground_endofpacket
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_valid;                                  // video_dual_clock_buffer_0:stream_out_valid -> video_vga_controller_0:valid
	wire  [29:0] video_dual_clock_buffer_0_avalon_dc_buffer_source_data;                                   // video_dual_clock_buffer_0:stream_out_data -> video_vga_controller_0:data
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_ready;                                  // video_vga_controller_0:ready -> video_dual_clock_buffer_0:stream_out_ready
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket;                          // video_dual_clock_buffer_0:stream_out_startofpacket -> video_vga_controller_0:startofpacket
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket;                            // video_dual_clock_buffer_0:stream_out_endofpacket -> video_vga_controller_0:endofpacket
	wire         video_pixel_buffer_dma_0_avalon_pixel_source_valid;                                       // video_pixel_buffer_dma_0:stream_valid -> video_rgb_resampler_0:stream_in_valid
	wire  [23:0] video_pixel_buffer_dma_0_avalon_pixel_source_data;                                        // video_pixel_buffer_dma_0:stream_data -> video_rgb_resampler_0:stream_in_data
	wire         video_pixel_buffer_dma_0_avalon_pixel_source_ready;                                       // video_rgb_resampler_0:stream_in_ready -> video_pixel_buffer_dma_0:stream_ready
	wire         video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket;                               // video_pixel_buffer_dma_0:stream_startofpacket -> video_rgb_resampler_0:stream_in_startofpacket
	wire         video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket;                                 // video_pixel_buffer_dma_0:stream_endofpacket -> video_rgb_resampler_0:stream_in_endofpacket
	wire         video_rgb_resampler_0_avalon_rgb_source_valid;                                            // video_rgb_resampler_0:stream_out_valid -> video_scaler_0:stream_in_valid
	wire  [29:0] video_rgb_resampler_0_avalon_rgb_source_data;                                             // video_rgb_resampler_0:stream_out_data -> video_scaler_0:stream_in_data
	wire         video_rgb_resampler_0_avalon_rgb_source_ready;                                            // video_scaler_0:stream_in_ready -> video_rgb_resampler_0:stream_out_ready
	wire         video_rgb_resampler_0_avalon_rgb_source_startofpacket;                                    // video_rgb_resampler_0:stream_out_startofpacket -> video_scaler_0:stream_in_startofpacket
	wire         video_rgb_resampler_0_avalon_rgb_source_endofpacket;                                      // video_rgb_resampler_0:stream_out_endofpacket -> video_scaler_0:stream_in_endofpacket
	wire         sys_sdram_pll_0_sys_clk_clk;                                                              // sys_sdram_pll_0:sys_clk_clk -> [irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:sys_sdram_pll_0_sys_clk_clk, nios2_gen2_0:clk, rst_controller:clk, rst_controller_001:clk]
	wire         video_pll_0_vga_clk_clk;                                                                  // video_pll_0:vga_clk_clk -> [rst_controller_004:clk, video_dual_clock_buffer_0:clk_stream_out, video_vga_controller_0:clk]
	wire         video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest;                             // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest -> video_pixel_buffer_dma_0:master_waitrequest
	wire  [31:0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata;                                // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata -> video_pixel_buffer_dma_0:master_readdata
	wire  [31:0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_address;                                 // video_pixel_buffer_dma_0:master_address -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_address
	wire         video_pixel_buffer_dma_0_avalon_pixel_dma_master_read;                                    // video_pixel_buffer_dma_0:master_read -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_read
	wire         video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid;                           // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid -> video_pixel_buffer_dma_0:master_readdatavalid
	wire         video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock;                                    // video_pixel_buffer_dma_0:master_arbiterlock -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock
	wire  [31:0] nios2_gen2_0_data_master_readdata;                                                        // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                                                     // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                                                     // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [28:0] nios2_gen2_0_data_master_address;                                                         // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                                                      // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                                            // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_readdatavalid;                                                   // mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire         nios2_gen2_0_data_master_write;                                                           // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                                                       // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                                                 // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                                              // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [28:0] nios2_gen2_0_instruction_master_address;                                                  // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                                                     // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;                                            // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire  [15:0] mm_interconnect_0_sram_0_avalon_sram_slave_readdata;                                      // sram_0:readdata -> mm_interconnect_0:sram_0_avalon_sram_slave_readdata
	wire  [19:0] mm_interconnect_0_sram_0_avalon_sram_slave_address;                                       // mm_interconnect_0:sram_0_avalon_sram_slave_address -> sram_0:address
	wire         mm_interconnect_0_sram_0_avalon_sram_slave_read;                                          // mm_interconnect_0:sram_0_avalon_sram_slave_read -> sram_0:read
	wire   [1:0] mm_interconnect_0_sram_0_avalon_sram_slave_byteenable;                                    // mm_interconnect_0:sram_0_avalon_sram_slave_byteenable -> sram_0:byteenable
	wire         mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid;                                 // sram_0:readdatavalid -> mm_interconnect_0:sram_0_avalon_sram_slave_readdatavalid
	wire         mm_interconnect_0_sram_0_avalon_sram_slave_write;                                         // mm_interconnect_0:sram_0_avalon_sram_slave_write -> sram_0:write
	wire  [15:0] mm_interconnect_0_sram_0_avalon_sram_slave_writedata;                                     // mm_interconnect_0:sram_0_avalon_sram_slave_writedata -> sram_0:writedata
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect;  // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect -> video_character_buffer_with_dma_0:buf_chipselect
	wire   [7:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata;    // video_character_buffer_with_dma_0:buf_readdata -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest; // video_character_buffer_with_dma_0:buf_waitrequest -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest
	wire  [12:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address;     // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_address -> video_character_buffer_with_dma_0:buf_address
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read;        // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_read -> video_character_buffer_with_dma_0:buf_read
	wire   [0:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable;  // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable -> video_character_buffer_with_dma_0:buf_byteenable
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write;       // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_write -> video_character_buffer_with_dma_0:buf_write
	wire   [7:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata;   // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata -> video_character_buffer_with_dma_0:buf_writedata
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect; // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect -> video_character_buffer_with_dma_0:ctrl_chipselect
	wire  [31:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata;   // video_character_buffer_with_dma_0:ctrl_readdata -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_readdata
	wire   [0:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address;    // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_address -> video_character_buffer_with_dma_0:ctrl_address
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read;       // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_read -> video_character_buffer_with_dma_0:ctrl_read
	wire   [3:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable; // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable -> video_character_buffer_with_dma_0:ctrl_byteenable
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write;      // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_write -> video_character_buffer_with_dma_0:ctrl_write
	wire  [31:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata;  // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_writedata -> video_character_buffer_with_dma_0:ctrl_writedata
	wire  [31:0] mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_readdata;                 // video_pixel_buffer_dma_0:slave_readdata -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_readdata
	wire   [1:0] mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_address;                  // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_address -> video_pixel_buffer_dma_0:slave_address
	wire         mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_read;                     // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_read -> video_pixel_buffer_dma_0:slave_read
	wire   [3:0] mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_byteenable;               // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_byteenable -> video_pixel_buffer_dma_0:slave_byteenable
	wire         mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_write;                    // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_write -> video_pixel_buffer_dma_0:slave_write
	wire  [31:0] mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_writedata;                // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_writedata -> video_pixel_buffer_dma_0:slave_writedata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;                               // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;                                 // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;                              // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;                                  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;                                     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;                                    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;                                // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_readdata;                        // video_rgb_resampler_0:slave_readdata -> mm_interconnect_0:video_rgb_resampler_0_avalon_rgb_slave_readdata
	wire         mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_read;                            // mm_interconnect_0:video_rgb_resampler_0_avalon_rgb_slave_read -> video_rgb_resampler_0:slave_read
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;                                  // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;                               // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;                               // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;                                   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;                                      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;                                // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;                                     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;                                 // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_sdram_controller_0_s1_chipselect;                                       // mm_interconnect_0:sdram_controller_0_s1_chipselect -> sdram_controller_0:az_cs
	wire  [31:0] mm_interconnect_0_sdram_controller_0_s1_readdata;                                         // sdram_controller_0:za_data -> mm_interconnect_0:sdram_controller_0_s1_readdata
	wire         mm_interconnect_0_sdram_controller_0_s1_waitrequest;                                      // sdram_controller_0:za_waitrequest -> mm_interconnect_0:sdram_controller_0_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_controller_0_s1_address;                                          // mm_interconnect_0:sdram_controller_0_s1_address -> sdram_controller_0:az_addr
	wire         mm_interconnect_0_sdram_controller_0_s1_read;                                             // mm_interconnect_0:sdram_controller_0_s1_read -> sdram_controller_0:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_controller_0_s1_byteenable;                                       // mm_interconnect_0:sdram_controller_0_s1_byteenable -> sdram_controller_0:az_be_n
	wire         mm_interconnect_0_sdram_controller_0_s1_readdatavalid;                                    // sdram_controller_0:za_valid -> mm_interconnect_0:sdram_controller_0_s1_readdatavalid
	wire         mm_interconnect_0_sdram_controller_0_s1_write;                                            // mm_interconnect_0:sdram_controller_0_s1_write -> sdram_controller_0:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_controller_0_s1_writedata;                                        // mm_interconnect_0:sdram_controller_0_s1_writedata -> sdram_controller_0:az_data
	wire         irq_mapper_receiver0_irq;                                                                 // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                                                     // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         video_scaler_0_avalon_scaler_source_valid;                                                // video_scaler_0:stream_out_valid -> avalon_st_adapter:in_0_valid
	wire  [29:0] video_scaler_0_avalon_scaler_source_data;                                                 // video_scaler_0:stream_out_data -> avalon_st_adapter:in_0_data
	wire         video_scaler_0_avalon_scaler_source_ready;                                                // avalon_st_adapter:in_0_ready -> video_scaler_0:stream_out_ready
	wire   [1:0] video_scaler_0_avalon_scaler_source_channel;                                              // video_scaler_0:stream_out_channel -> avalon_st_adapter:in_0_channel
	wire         video_scaler_0_avalon_scaler_source_startofpacket;                                        // video_scaler_0:stream_out_startofpacket -> avalon_st_adapter:in_0_startofpacket
	wire         video_scaler_0_avalon_scaler_source_endofpacket;                                          // video_scaler_0:stream_out_endofpacket -> avalon_st_adapter:in_0_endofpacket
	wire         avalon_st_adapter_out_0_valid;                                                            // avalon_st_adapter:out_0_valid -> video_alpha_blender_0:background_valid
	wire  [29:0] avalon_st_adapter_out_0_data;                                                             // avalon_st_adapter:out_0_data -> video_alpha_blender_0:background_data
	wire         avalon_st_adapter_out_0_ready;                                                            // video_alpha_blender_0:background_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                                                    // avalon_st_adapter:out_0_startofpacket -> video_alpha_blender_0:background_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                                                      // avalon_st_adapter:out_0_endofpacket -> video_alpha_blender_0:background_endofpacket
	wire         rst_controller_reset_out_reset;                                                           // rst_controller:reset_out -> [jtag_uart_0:rst_n, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                                                       // rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                                                   // rst_controller_001:reset_req -> [nios2_gen2_0:reset_req, rst_translator:reset_req_in]
	wire         sys_sdram_pll_0_reset_source_reset;                                                       // sys_sdram_pll_0:reset_source_reset -> rst_controller_001:reset_in0
	wire         rst_controller_002_reset_out_reset;                                                       // rst_controller_002:reset_out -> [mm_interconnect_0:sdram_controller_0_reset_reset_bridge_in_reset_reset, sdram_controller_0:reset_n]
	wire         rst_controller_003_reset_out_reset;                                                       // rst_controller_003:reset_out -> [avalon_st_adapter:in_rst_0_reset, mm_interconnect_0:video_pixel_buffer_dma_0_reset_reset_bridge_in_reset_reset, sram_0:reset, sys_sdram_pll_0:ref_reset_reset, video_alpha_blender_0:reset, video_character_buffer_with_dma_0:reset, video_dual_clock_buffer_0:reset_stream_in, video_pixel_buffer_dma_0:reset, video_pll_0:ref_reset_reset, video_rgb_resampler_0:reset, video_scaler_0:reset]
	wire         rst_controller_004_reset_out_reset;                                                       // rst_controller_004:reset_out -> [video_dual_clock_buffer_0:reset_stream_out, video_vga_controller_0:reset]
	wire         video_pll_0_reset_source_reset;                                                           // video_pll_0:reset_source_reset -> rst_controller_004:reset_in0

	nios_system_jtag_uart_0 jtag_uart_0 (
		.clk            (sys_sdram_pll_0_sys_clk_clk),                                 //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	nios_system_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (sys_sdram_pll_0_sys_clk_clk),                                //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	nios_system_sdram_controller_0 sdram_controller_0 (
		.clk            (sdram_clk_clk),                                         //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),                   // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controller_0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controller_0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controller_0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controller_0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controller_0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controller_0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controller_0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controller_0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controller_0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (new_sdram_controller_0_wire_addr),                      //  wire.export
		.zs_ba          (new_sdram_controller_0_wire_ba),                        //      .export
		.zs_cas_n       (new_sdram_controller_0_wire_cas_n),                     //      .export
		.zs_cke         (new_sdram_controller_0_wire_cke),                       //      .export
		.zs_cs_n        (new_sdram_controller_0_wire_cs_n),                      //      .export
		.zs_dq          (new_sdram_controller_0_wire_dq),                        //      .export
		.zs_dqm         (new_sdram_controller_0_wire_dqm),                       //      .export
		.zs_ras_n       (new_sdram_controller_0_wire_ras_n),                     //      .export
		.zs_we_n        (new_sdram_controller_0_wire_we_n)                       //      .export
	);

	nios_system_sram_0 sram_0 (
		.clk           (clk_clk),                                                  //                clk.clk
		.reset         (rst_controller_003_reset_out_reset),                       //              reset.reset
		.SRAM_DQ       (sram_DQ),                                                  // external_interface.export
		.SRAM_ADDR     (sram_ADDR),                                                //                   .export
		.SRAM_LB_N     (sram_LB_N),                                                //                   .export
		.SRAM_UB_N     (sram_UB_N),                                                //                   .export
		.SRAM_CE_N     (sram_CE_N),                                                //                   .export
		.SRAM_OE_N     (sram_OE_N),                                                //                   .export
		.SRAM_WE_N     (sram_WE_N),                                                //                   .export
		.address       (mm_interconnect_0_sram_0_avalon_sram_slave_address),       //  avalon_sram_slave.address
		.byteenable    (mm_interconnect_0_sram_0_avalon_sram_slave_byteenable),    //                   .byteenable
		.read          (mm_interconnect_0_sram_0_avalon_sram_slave_read),          //                   .read
		.write         (mm_interconnect_0_sram_0_avalon_sram_slave_write),         //                   .write
		.writedata     (mm_interconnect_0_sram_0_avalon_sram_slave_writedata),     //                   .writedata
		.readdata      (mm_interconnect_0_sram_0_avalon_sram_slave_readdata),      //                   .readdata
		.readdatavalid (mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid)  //                   .readdatavalid
	);

	nios_system_sys_sdram_pll_0 sys_sdram_pll_0 (
		.ref_clk_clk        (clk_clk),                            //      ref_clk.clk
		.ref_reset_reset    (rst_controller_003_reset_out_reset), //    ref_reset.reset
		.sys_clk_clk        (sys_sdram_pll_0_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                      //    sdram_clk.clk
		.reset_source_reset (sys_sdram_pll_0_reset_source_reset)  // reset_source.reset
	);

	nios_system_video_alpha_blender_0 video_alpha_blender_0 (
		.clk                      (clk_clk),                                                            //                    clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                 //                  reset.reset
		.foreground_data          (video_character_buffer_with_dma_0_avalon_char_source_data),          // avalon_foreground_sink.data
		.foreground_startofpacket (video_character_buffer_with_dma_0_avalon_char_source_startofpacket), //                       .startofpacket
		.foreground_endofpacket   (video_character_buffer_with_dma_0_avalon_char_source_endofpacket),   //                       .endofpacket
		.foreground_valid         (video_character_buffer_with_dma_0_avalon_char_source_valid),         //                       .valid
		.foreground_ready         (video_character_buffer_with_dma_0_avalon_char_source_ready),         //                       .ready
		.background_data          (avalon_st_adapter_out_0_data),                                       // avalon_background_sink.data
		.background_startofpacket (avalon_st_adapter_out_0_startofpacket),                              //                       .startofpacket
		.background_endofpacket   (avalon_st_adapter_out_0_endofpacket),                                //                       .endofpacket
		.background_valid         (avalon_st_adapter_out_0_valid),                                      //                       .valid
		.background_ready         (avalon_st_adapter_out_0_ready),                                      //                       .ready
		.output_ready             (video_alpha_blender_0_avalon_blended_source_ready),                  //  avalon_blended_source.ready
		.output_data              (video_alpha_blender_0_avalon_blended_source_data),                   //                       .data
		.output_startofpacket     (video_alpha_blender_0_avalon_blended_source_startofpacket),          //                       .startofpacket
		.output_endofpacket       (video_alpha_blender_0_avalon_blended_source_endofpacket),            //                       .endofpacket
		.output_valid             (video_alpha_blender_0_avalon_blended_source_valid)                   //                       .valid
	);

	nios_system_video_character_buffer_with_dma_0 video_character_buffer_with_dma_0 (
		.clk                  (clk_clk),                                                                                  //                       clk.clk
		.reset                (rst_controller_003_reset_out_reset),                                                       //                     reset.reset
		.ctrl_address         (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address),    // avalon_char_control_slave.address
		.ctrl_byteenable      (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable), //                          .byteenable
		.ctrl_chipselect      (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect), //                          .chipselect
		.ctrl_read            (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read),       //                          .read
		.ctrl_write           (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write),      //                          .write
		.ctrl_writedata       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata),  //                          .writedata
		.ctrl_readdata        (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata),   //                          .readdata
		.buf_byteenable       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable),  //  avalon_char_buffer_slave.byteenable
		.buf_chipselect       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect),  //                          .chipselect
		.buf_read             (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read),        //                          .read
		.buf_write            (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write),       //                          .write
		.buf_writedata        (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata),   //                          .writedata
		.buf_readdata         (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata),    //                          .readdata
		.buf_waitrequest      (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest), //                          .waitrequest
		.buf_address          (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address),     //                          .address
		.stream_ready         (video_character_buffer_with_dma_0_avalon_char_source_ready),                               //        avalon_char_source.ready
		.stream_startofpacket (video_character_buffer_with_dma_0_avalon_char_source_startofpacket),                       //                          .startofpacket
		.stream_endofpacket   (video_character_buffer_with_dma_0_avalon_char_source_endofpacket),                         //                          .endofpacket
		.stream_valid         (video_character_buffer_with_dma_0_avalon_char_source_valid),                               //                          .valid
		.stream_data          (video_character_buffer_with_dma_0_avalon_char_source_data)                                 //                          .data
	);

	nios_system_video_dual_clock_buffer_0 video_dual_clock_buffer_0 (
		.clk_stream_in            (clk_clk),                                                         //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_003_reset_out_reset),                              //         reset_stream_in.reset
		.clk_stream_out           (video_pll_0_vga_clk_clk),                                         //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_004_reset_out_reset),                              //        reset_stream_out.reset
		.stream_in_ready          (video_alpha_blender_0_avalon_blended_source_ready),               //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (video_alpha_blender_0_avalon_blended_source_startofpacket),       //                        .startofpacket
		.stream_in_endofpacket    (video_alpha_blender_0_avalon_blended_source_endofpacket),         //                        .endofpacket
		.stream_in_valid          (video_alpha_blender_0_avalon_blended_source_valid),               //                        .valid
		.stream_in_data           (video_alpha_blender_0_avalon_blended_source_data),                //                        .data
		.stream_out_ready         (video_dual_clock_buffer_0_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (video_dual_clock_buffer_0_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (video_dual_clock_buffer_0_avalon_dc_buffer_source_data)           //                        .data
	);

	nios_system_video_pixel_buffer_dma_0 video_pixel_buffer_dma_0 (
		.clk                  (clk_clk),                                                                    //                     clk.clk
		.reset                (rst_controller_003_reset_out_reset),                                         //                   reset.reset
		.master_readdatavalid (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid),             // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest),               //                        .waitrequest
		.master_address       (video_pixel_buffer_dma_0_avalon_pixel_dma_master_address),                   //                        .address
		.master_arbiterlock   (video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock),                      //                        .lock
		.master_read          (video_pixel_buffer_dma_0_avalon_pixel_dma_master_read),                      //                        .read
		.master_readdata      (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata),                  //                        .readdata
		.slave_address        (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_address),    //    avalon_control_slave.address
		.slave_byteenable     (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_byteenable), //                        .byteenable
		.slave_read           (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_read),       //                        .read
		.slave_write          (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_write),      //                        .write
		.slave_writedata      (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_writedata),  //                        .writedata
		.slave_readdata       (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_readdata),   //                        .readdata
		.stream_ready         (video_pixel_buffer_dma_0_avalon_pixel_source_ready),                         //     avalon_pixel_source.ready
		.stream_startofpacket (video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket),                 //                        .startofpacket
		.stream_endofpacket   (video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket),                   //                        .endofpacket
		.stream_valid         (video_pixel_buffer_dma_0_avalon_pixel_source_valid),                         //                        .valid
		.stream_data          (video_pixel_buffer_dma_0_avalon_pixel_source_data)                           //                        .data
	);

	nios_system_video_pll_0 video_pll_0 (
		.ref_clk_clk        (clk_clk),                            //      ref_clk.clk
		.ref_reset_reset    (rst_controller_003_reset_out_reset), //    ref_reset.reset
		.video_in_clk_clk   (),                                   // video_in_clk.clk
		.vga_clk_clk        (video_pll_0_vga_clk_clk),            //      vga_clk.clk
		.lcd_clk_clk        (),                                   //      lcd_clk.clk
		.reset_source_reset (video_pll_0_reset_source_reset)      // reset_source.reset
	);

	nios_system_video_rgb_resampler_0 video_rgb_resampler_0 (
		.clk                      (clk_clk),                                                           //               clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                //             reset.reset
		.stream_in_startofpacket  (video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket),        //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket),          //                  .endofpacket
		.stream_in_valid          (video_pixel_buffer_dma_0_avalon_pixel_source_valid),                //                  .valid
		.stream_in_ready          (video_pixel_buffer_dma_0_avalon_pixel_source_ready),                //                  .ready
		.stream_in_data           (video_pixel_buffer_dma_0_avalon_pixel_source_data),                 //                  .data
		.slave_read               (mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_read),     //  avalon_rgb_slave.read
		.slave_readdata           (mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_readdata), //                  .readdata
		.stream_out_ready         (video_rgb_resampler_0_avalon_rgb_source_ready),                     // avalon_rgb_source.ready
		.stream_out_startofpacket (video_rgb_resampler_0_avalon_rgb_source_startofpacket),             //                  .startofpacket
		.stream_out_endofpacket   (video_rgb_resampler_0_avalon_rgb_source_endofpacket),               //                  .endofpacket
		.stream_out_valid         (video_rgb_resampler_0_avalon_rgb_source_valid),                     //                  .valid
		.stream_out_data          (video_rgb_resampler_0_avalon_rgb_source_data)                       //                  .data
	);

	nios_system_video_scaler_0 video_scaler_0 (
		.clk                      (clk_clk),                                               //                  clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                    //                reset.reset
		.stream_in_startofpacket  (video_rgb_resampler_0_avalon_rgb_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (video_rgb_resampler_0_avalon_rgb_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (video_rgb_resampler_0_avalon_rgb_source_valid),         //                     .valid
		.stream_in_ready          (video_rgb_resampler_0_avalon_rgb_source_ready),         //                     .ready
		.stream_in_data           (video_rgb_resampler_0_avalon_rgb_source_data),          //                     .data
		.stream_out_ready         (video_scaler_0_avalon_scaler_source_ready),             // avalon_scaler_source.ready
		.stream_out_startofpacket (video_scaler_0_avalon_scaler_source_startofpacket),     //                     .startofpacket
		.stream_out_endofpacket   (video_scaler_0_avalon_scaler_source_endofpacket),       //                     .endofpacket
		.stream_out_valid         (video_scaler_0_avalon_scaler_source_valid),             //                     .valid
		.stream_out_data          (video_scaler_0_avalon_scaler_source_data),              //                     .data
		.stream_out_channel       (video_scaler_0_avalon_scaler_source_channel)            //                     .channel
	);

	nios_system_video_vga_controller_0 video_vga_controller_0 (
		.clk           (video_pll_0_vga_clk_clk),                                         //                clk.clk
		.reset         (rst_controller_004_reset_out_reset),                              //              reset.reset
		.data          (video_dual_clock_buffer_0_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (video_dual_clock_buffer_0_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (video_dual_clock_buffer_0_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_CLK),                                                         // external_interface.export
		.VGA_HS        (vga_HS),                                                          //                   .export
		.VGA_VS        (vga_VS),                                                          //                   .export
		.VGA_BLANK     (vga_BLANK),                                                       //                   .export
		.VGA_SYNC      (vga_SYNC),                                                        //                   .export
		.VGA_R         (vga_R),                                                           //                   .export
		.VGA_G         (vga_G),                                                           //                   .export
		.VGA_B         (vga_B)                                                            //                   .export
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                                          (clk_clk),                                                                                  //                                                   clk_0_clk.clk
		.sys_sdram_pll_0_sdram_clk_clk                                          (sdram_clk_clk),                                                                            //                                   sys_sdram_pll_0_sdram_clk.clk
		.sys_sdram_pll_0_sys_clk_clk                                            (sys_sdram_pll_0_sys_clk_clk),                                                              //                                     sys_sdram_pll_0_sys_clk.clk
		.jtag_uart_0_reset_reset_bridge_in_reset_reset                          (rst_controller_reset_out_reset),                                                           //                     jtag_uart_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset                         (rst_controller_001_reset_out_reset),                                                       //                    nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.sdram_controller_0_reset_reset_bridge_in_reset_reset                   (rst_controller_002_reset_out_reset),                                                       //              sdram_controller_0_reset_reset_bridge_in_reset.reset
		.video_pixel_buffer_dma_0_reset_reset_bridge_in_reset_reset             (rst_controller_003_reset_out_reset),                                                       //        video_pixel_buffer_dma_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                                       (nios2_gen2_0_data_master_address),                                                         //                                    nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                                   (nios2_gen2_0_data_master_waitrequest),                                                     //                                                            .waitrequest
		.nios2_gen2_0_data_master_byteenable                                    (nios2_gen2_0_data_master_byteenable),                                                      //                                                            .byteenable
		.nios2_gen2_0_data_master_read                                          (nios2_gen2_0_data_master_read),                                                            //                                                            .read
		.nios2_gen2_0_data_master_readdata                                      (nios2_gen2_0_data_master_readdata),                                                        //                                                            .readdata
		.nios2_gen2_0_data_master_readdatavalid                                 (nios2_gen2_0_data_master_readdatavalid),                                                   //                                                            .readdatavalid
		.nios2_gen2_0_data_master_write                                         (nios2_gen2_0_data_master_write),                                                           //                                                            .write
		.nios2_gen2_0_data_master_writedata                                     (nios2_gen2_0_data_master_writedata),                                                       //                                                            .writedata
		.nios2_gen2_0_data_master_debugaccess                                   (nios2_gen2_0_data_master_debugaccess),                                                     //                                                            .debugaccess
		.nios2_gen2_0_instruction_master_address                                (nios2_gen2_0_instruction_master_address),                                                  //                             nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest                            (nios2_gen2_0_instruction_master_waitrequest),                                              //                                                            .waitrequest
		.nios2_gen2_0_instruction_master_read                                   (nios2_gen2_0_instruction_master_read),                                                     //                                                            .read
		.nios2_gen2_0_instruction_master_readdata                               (nios2_gen2_0_instruction_master_readdata),                                                 //                                                            .readdata
		.nios2_gen2_0_instruction_master_readdatavalid                          (nios2_gen2_0_instruction_master_readdatavalid),                                            //                                                            .readdatavalid
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_address               (video_pixel_buffer_dma_0_avalon_pixel_dma_master_address),                                 //            video_pixel_buffer_dma_0_avalon_pixel_dma_master.address
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest           (video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest),                             //                                                            .waitrequest
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_read                  (video_pixel_buffer_dma_0_avalon_pixel_dma_master_read),                                    //                                                            .read
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata              (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata),                                //                                                            .readdata
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid         (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid),                           //                                                            .readdatavalid
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock                  (video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock),                                    //                                                            .lock
		.jtag_uart_0_avalon_jtag_slave_address                                  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),                                  //                               jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                                    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),                                    //                                                            .write
		.jtag_uart_0_avalon_jtag_slave_read                                     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),                                     //                                                            .read
		.jtag_uart_0_avalon_jtag_slave_readdata                                 (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),                                 //                                                            .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                                (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),                                //                                                            .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),                              //                                                            .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),                               //                                                            .chipselect
		.nios2_gen2_0_debug_mem_slave_address                                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),                                   //                                nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                                     (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),                                     //                                                            .write
		.nios2_gen2_0_debug_mem_slave_read                                      (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),                                      //                                                            .read
		.nios2_gen2_0_debug_mem_slave_readdata                                  (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),                                  //                                                            .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                                 (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),                                 //                                                            .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable                                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),                                //                                                            .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest                               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),                               //                                                            .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess                               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),                               //                                                            .debugaccess
		.sdram_controller_0_s1_address                                          (mm_interconnect_0_sdram_controller_0_s1_address),                                          //                                       sdram_controller_0_s1.address
		.sdram_controller_0_s1_write                                            (mm_interconnect_0_sdram_controller_0_s1_write),                                            //                                                            .write
		.sdram_controller_0_s1_read                                             (mm_interconnect_0_sdram_controller_0_s1_read),                                             //                                                            .read
		.sdram_controller_0_s1_readdata                                         (mm_interconnect_0_sdram_controller_0_s1_readdata),                                         //                                                            .readdata
		.sdram_controller_0_s1_writedata                                        (mm_interconnect_0_sdram_controller_0_s1_writedata),                                        //                                                            .writedata
		.sdram_controller_0_s1_byteenable                                       (mm_interconnect_0_sdram_controller_0_s1_byteenable),                                       //                                                            .byteenable
		.sdram_controller_0_s1_readdatavalid                                    (mm_interconnect_0_sdram_controller_0_s1_readdatavalid),                                    //                                                            .readdatavalid
		.sdram_controller_0_s1_waitrequest                                      (mm_interconnect_0_sdram_controller_0_s1_waitrequest),                                      //                                                            .waitrequest
		.sdram_controller_0_s1_chipselect                                       (mm_interconnect_0_sdram_controller_0_s1_chipselect),                                       //                                                            .chipselect
		.sram_0_avalon_sram_slave_address                                       (mm_interconnect_0_sram_0_avalon_sram_slave_address),                                       //                                    sram_0_avalon_sram_slave.address
		.sram_0_avalon_sram_slave_write                                         (mm_interconnect_0_sram_0_avalon_sram_slave_write),                                         //                                                            .write
		.sram_0_avalon_sram_slave_read                                          (mm_interconnect_0_sram_0_avalon_sram_slave_read),                                          //                                                            .read
		.sram_0_avalon_sram_slave_readdata                                      (mm_interconnect_0_sram_0_avalon_sram_slave_readdata),                                      //                                                            .readdata
		.sram_0_avalon_sram_slave_writedata                                     (mm_interconnect_0_sram_0_avalon_sram_slave_writedata),                                     //                                                            .writedata
		.sram_0_avalon_sram_slave_byteenable                                    (mm_interconnect_0_sram_0_avalon_sram_slave_byteenable),                                    //                                                            .byteenable
		.sram_0_avalon_sram_slave_readdatavalid                                 (mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid),                                 //                                                            .readdatavalid
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_address     (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address),     //  video_character_buffer_with_dma_0_avalon_char_buffer_slave.address
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_write       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write),       //                                                            .write
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_read        (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read),        //                                                            .read
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata    (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata),    //                                                            .readdata
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata   (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata),   //                                                            .writedata
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable  (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable),  //                                                            .byteenable
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest), //                                                            .waitrequest
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect  (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect),  //                                                            .chipselect
		.video_character_buffer_with_dma_0_avalon_char_control_slave_address    (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address),    // video_character_buffer_with_dma_0_avalon_char_control_slave.address
		.video_character_buffer_with_dma_0_avalon_char_control_slave_write      (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write),      //                                                            .write
		.video_character_buffer_with_dma_0_avalon_char_control_slave_read       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read),       //                                                            .read
		.video_character_buffer_with_dma_0_avalon_char_control_slave_readdata   (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata),   //                                                            .readdata
		.video_character_buffer_with_dma_0_avalon_char_control_slave_writedata  (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata),  //                                                            .writedata
		.video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable), //                                                            .byteenable
		.video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect), //                                                            .chipselect
		.video_pixel_buffer_dma_0_avalon_control_slave_address                  (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_address),                  //               video_pixel_buffer_dma_0_avalon_control_slave.address
		.video_pixel_buffer_dma_0_avalon_control_slave_write                    (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_write),                    //                                                            .write
		.video_pixel_buffer_dma_0_avalon_control_slave_read                     (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_read),                     //                                                            .read
		.video_pixel_buffer_dma_0_avalon_control_slave_readdata                 (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_readdata),                 //                                                            .readdata
		.video_pixel_buffer_dma_0_avalon_control_slave_writedata                (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_writedata),                //                                                            .writedata
		.video_pixel_buffer_dma_0_avalon_control_slave_byteenable               (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_byteenable),               //                                                            .byteenable
		.video_rgb_resampler_0_avalon_rgb_slave_read                            (mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_read),                            //                      video_rgb_resampler_0_avalon_rgb_slave.read
		.video_rgb_resampler_0_avalon_rgb_slave_readdata                        (mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_readdata)                         //                                                            .readdata
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (sys_sdram_pll_0_sys_clk_clk),        //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	nios_system_avalon_st_adapter #(
		.inBitsPerSymbol (10),
		.inUsePackets    (1),
		.inDataWidth     (30),
		.inChannelWidth  (2),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (30),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (clk_clk),                                           // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_003_reset_out_reset),                // in_rst_0.reset
		.in_0_data           (video_scaler_0_avalon_scaler_source_data),          //     in_0.data
		.in_0_valid          (video_scaler_0_avalon_scaler_source_valid),         //         .valid
		.in_0_ready          (video_scaler_0_avalon_scaler_source_ready),         //         .ready
		.in_0_startofpacket  (video_scaler_0_avalon_scaler_source_startofpacket), //         .startofpacket
		.in_0_endofpacket    (video_scaler_0_avalon_scaler_source_endofpacket),   //         .endofpacket
		.in_0_channel        (video_scaler_0_avalon_scaler_source_channel),       //         .channel
		.out_0_data          (avalon_st_adapter_out_0_data),                      //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),                     //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),                     //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket),             //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket)                //         .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (sys_sdram_pll_0_sys_clk_clk),    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (sys_sdram_pll_0_reset_source_reset),     // reset_in0.reset
		.clk            (sys_sdram_pll_0_sys_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (sdram_clk_clk),                      //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (video_pll_0_reset_source_reset),     // reset_in0.reset
		.clk            (video_pll_0_vga_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
